module shifts;
reg signed [7:0]a;

initial
begin
	a=8'b1101_0011;
	$display("logical left shift=%b",a<<1);
	$display("logical right shift=%b",a>>1);
	$display("arithmatic left shift=%b",a<<<1);
	$display("arithmatic right shift=%b",a>>>1);

	a=8'b0101_0011;
	$display("logical left shift=%b",a<<1);
	$display("logical right shift=%b",a>>1);
	$display("arithmatic left shift=%b",a<<<1);
	$display("arithmatic right shift=%b",a>>>1);

	a=8'b1101_0010;
	$display("logical left shift=%b",a<<1);
	$display("logical right shift=%b",a>>1);
	$display("arithmatic left shift=%b",a<<<1);
	$display("arithmatic right shift=%b",a>>>1);

	a=8'b0101_0010;
	$display("logical left shift=%b",a<<1);
	$display("logical right shift=%b",a>>1);
	$display("arithmatic left shift=%b",a<<<1);
	$display("arithmatic right shift=%b",a>>>1);
end 
endmodule
