module b2gdataflow(bin, gray);
	/////////// 
endmodule
